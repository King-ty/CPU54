`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/05/29 12:25:58
// Design Name: 
// Module Name: IMEM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module IMEM(
    input [10:0] addr,	//ָ���ַ
    output [31:0] instr	//ָ������
    );

    // reg [31:0] temp;//?

    IMEM_ROM I_ROM (
        .a(addr),      // input wire [10 : 0] a
        .spo(instr)  // output wire [31 : 0] spo
    );
endmodule
